library verilog;
use verilog.vl_types.all;
entity ex04 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        F               : out    vl_logic
    );
end ex04;
