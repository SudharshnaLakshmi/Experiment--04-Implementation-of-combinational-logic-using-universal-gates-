library verilog;
use verilog.vl_types.all;
entity ex04_vlg_vec_tst is
end ex04_vlg_vec_tst;
